module HDSimulado
#(parameter DATA_WIDTH=32, parameter ADDR_WIDTH=9)
(
	input [(DATA_WIDTH-1):0] data,
	input [(ADDR_WIDTH-1):0] addr,
	input we, clk,
	output [(DATA_WIDTH-1):0] q
);

	// Declare the RAM variable
	reg [DATA_WIDTH-1:0] HardDisk[2**ADDR_WIDTH-1:0];

	// Variable to hold the registered read address
	reg [ADDR_WIDTH-1:0] addr_reg;

	initial 
	begin : INIT
		integer i;
		HardDisk[ 0] = 32'B01011100000000000000000000000000; // HD_HEAD
		HardDisk[ 1] = 32'B01010100000000000000000000000000; // BEGIN_FILE
		HardDisk[ 2] = 32'B00001000000000010000000000000100; // addi	$ra $zero 4
		HardDisk[ 3] = 32'B00001000000111110000000000110110; // addi	$sp $zero 54
		HardDisk[ 4] = 32'B00010100000000000000000000000011; // jump	main
		HardDisk[ 5] = 32'B00110000000000000000000000000000; // nop	main
		HardDisk[ 6] = 32'B00001000000010000000000000000110; // addi	$t0 $zero 6
		HardDisk[ 7] = 32'B00011100000010000000000000000001; // sw	$t0 1($zero)
		HardDisk[ 8] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		HardDisk[ 9] = 32'B00011100000010000000000000000000; // sw	$t0 0($zero)
		HardDisk[10] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		HardDisk[11] = 32'B00011100000010000000000000000010; // sw	$t0 2($zero)
		HardDisk[12] = 32'B00110000000000000000000000000000; // nop	L0
		HardDisk[13] = 32'B00011000000101000000000000000000; // lw	$s0 0($zero)
		HardDisk[14] = 32'B00011000000101010000000000000001; // lw	$s1 1($zero)
		HardDisk[15] = 32'B00010010100101010100000000000000; // slt	$t0 $s0 $s1
		HardDisk[16] = 32'B00101001000000000000000000011101; // beq	$t0 0 L1
		HardDisk[17] = 32'B00001000000010010000000000000010; // addi	$t1 $zero 2
		HardDisk[18] = 32'B00011000000101010000000000000010; // lw	$s1 2($zero)
		HardDisk[19] = 32'B00000001001101010101000000000010; // mult	$t2 $t1 $s1
		HardDisk[20] = 32'B00011100000010100000000000000010; // sw	$t2 2($zero)
		HardDisk[21] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		HardDisk[22] = 32'B00011000000101000000000000000000; // lw	$s0 0($zero)
		HardDisk[23] = 32'B00000001000101000100100000000000; // add	$t1 $s0 $t0
		HardDisk[24] = 32'B00011100000010010000000000000000; // sw	$t1 0($zero)
		HardDisk[25] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		HardDisk[26] = 32'B00011000000101000000000000000010; // lw	$s0 2($zero)
		HardDisk[27] = 32'B00000010100010000100100000000001; // sub	$t1 $s0 $t0
		HardDisk[28] = 32'B00001101001000100000000000000000; // move	$a0 $t1 
		HardDisk[29] = 32'B00100100010000000000000000000000; // out	$a0  
		HardDisk[30] = 32'B00010100000000000000000000001010; // jump	L0
		HardDisk[31] = 32'B00110000000000000000000000000000; // nop	L1
		HardDisk[32] = 32'B00010100000000000000000000011110; // halt	  
		HardDisk[33] = 32'B01011000000000000000000000000000; // END_FILE
		HardDisk[34] = 32'B01100000000000000000000000000000; // HD_END
	end 

	always @ (posedge clk)
	begin
	
		// Write
		if (we)
			HardDisk[addr] <= data;

		addr_reg <= addr;
	end
 
	assign q = HardDisk[addr_reg];

endmodule
