module ShiftLeft2(Imediato,Output);
	input[31:0] Imediato;
	output reg[31:0] Output;
endmodule




