module ControleULA(OpALU,OpCode,funct);
	input [3:0] OpALU;
	output reg [5:0] OpCode,funct;



endmodule
