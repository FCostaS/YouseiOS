module HDSimulado
#(parameter DATA_WIDTH=32, parameter ADDR_WIDTH=9)
(
	input [(DATA_WIDTH-1):0] data,
	input [(ADDR_WIDTH-1):0] addr,
	input we, clk,
	output [(DATA_WIDTH-1):0] q
);

	// Declare the RAM variable
	reg [DATA_WIDTH-1:0] ram[2**ADDR_WIDTH-1:0];

	// Variable to hold the registered read address
	reg [ADDR_WIDTH-1:0] addr_reg;

	initial 
	begin : INIT
		integer i;
		ram[ 0] = 32'B01010100000000000000000000000000; // begin file	  
		ram[ 1] = 32'B00001000000000010000000000001000; // addi	$ra $zero 8
		ram[ 2] = 32'B00001000000111110000000000111010; // addi	$sp $zero 58
		ram[ 3] = 32'B00010100000000000000000000101001; // jump	main
		ram[ 4] = 32'B00110000000000000000000000000000; // nop	Combinatoria
		ram[ 5] = 32'B00011100000000100000000000000000; // sw	$a0 0($zero)
		ram[ 6] = 32'B00011100000000110000000000000001; // sw	$a1 1($zero)
		ram[ 7] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[ 8] = 32'B00011100000010000000000000000010; // sw	$t0 2($zero)
		ram[ 9] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[10] = 32'B00011100000010000000000000000011; // sw	$t0 3($zero)
		ram[11] = 32'B00110000000000000000000000000000; // nop	L0
		ram[12] = 32'B00001000000010000000000000000000; // addi	$t0 $zero 0
		ram[13] = 32'B00011000000101000000000000000001; // lw	$s0 1($zero)
		ram[14] = 32'B00111110100010000100100000000000; // sbt	$t1 $s0 $t0
		ram[15] = 32'B00101001001000000000000000100001; // beq	$t1 0 L1
		ram[16] = 32'B00011000000101000000000000000010; // lw	$s0 2($zero)
		ram[17] = 32'B00011000000101010000000000000000; // lw	$s1 0($zero)
		ram[18] = 32'B00000010100101010101000000000010; // mult	$t2 $s0 $s1
		ram[19] = 32'B00011100000010100000000000000010; // sw	$t2 2($zero)
		ram[20] = 32'B00011000000101000000000000000011; // lw	$s0 3($zero)
		ram[21] = 32'B00011000000101010000000000000001; // lw	$s1 1($zero)
		ram[22] = 32'B00000010100101010100000000000010; // mult	$t0 $s0 $s1
		ram[23] = 32'B00011100000010000000000000000011; // sw	$t0 3($zero)
		ram[24] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[25] = 32'B00011000000101000000000000000000; // lw	$s0 0($zero)
		ram[26] = 32'B00000010100010000100100000000001; // sub	$t1 $s0 $t0
		ram[27] = 32'B00011100000010010000000000000000; // sw	$t1 0($zero)
		ram[28] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[29] = 32'B00011000000101000000000000000001; // lw	$s0 1($zero)
		ram[30] = 32'B00000010100010000100100000000001; // sub	$t1 $s0 $t0
		ram[31] = 32'B00011100000010010000000000000001; // sw	$t1 1($zero)
		ram[32] = 32'B00010100000000000000000000001011; // jump	L0
		ram[33] = 32'B00110000000000000000000000000000; // nop	L1
		ram[34] = 32'B00011000000101000000000000000010; // lw	$s0 2($zero)
		ram[35] = 32'B00011000000101010000000000000011; // lw	$s1 3($zero)
		ram[36] = 32'B00000010100101010100000000000011; // div	$t0 $s0 $s1
		ram[37] = 32'B00001101000111100000000000000000; // move	$v0 $t0 
		ram[38] = 32'B01010000001000010000000000000001; // subi	$ra $ra 1
		ram[39] = 32'B00011000001101000000000000000000; // lw	$s0 0($ra)
		ram[40] = 32'B01001110100000000000000000000000; // jr	$s0  
		ram[41] = 32'B00110000000000000000000000000000; // nop	main
		ram[42] = 32'B00001000000010010000000000001111; // addi	$t1 $zero 15
		ram[43] = 32'B00011100000010010000000000000100; // sw	$t1 4($zero)
		ram[44] = 32'B00001000000010000000000000000110; // addi	$t0 $zero 6
		ram[45] = 32'B00011100000010000000000000000101; // sw	$t0 5($zero)
		ram[46] = 32'B00011000000101010000000000000100; // lw	$s1 4($zero)
		ram[47] = 32'B00001110101000100000000000000000; // move	$a0 $s1 
		ram[48] = 32'B00011000000101010000000000000101; // lw	$s1 5($zero)
		ram[49] = 32'B00001110101000110000000000000000; // move	$a1 $s1 
		ram[50] = 32'B00001000000101000000000000110110; // addi	$s0 $zero 54
		ram[51] = 32'B00011100001101000000000000000000; // sw	$s0 0($ra)
		ram[52] = 32'B00001000001000010000000000000001; // addi	$ra $ra 1
		ram[53] = 32'B00010100000000000000000000000100; // jump	Combinatoria
		ram[54] = 32'B00001111110001000000000000000000; // move	$a2 $v0 
		ram[55] = 32'B00100100100000000000000000000000; // out	$a2   
		ram[56] = 32'B01110000000000000000000000000001; // Set PID 1	  
		ram[57] = 32'B01011000000000000000000000111001; // end file
		ram[58] = 32'B01010100000000000000000000000000; // begin file	  
		ram[59] = 32'B00001000000000010000000000000100; // addi	$ra $zero 4
		ram[60] = 32'B00001000000111110000000000110110; // addi	$sp $zero 54
		ram[61] = 32'B00010100000000000000000000000100; // jump	main
		ram[62] = 32'B00110000000000000000000000000000; // nop	main
		ram[63] = 32'B00001000000010000000000000010100; // addi	$t0 $zero 20
		ram[64] = 32'B00011100000010000000000000000000; // sw	$t0 0($zero)
		ram[65] = 32'B00001000000010000000000001000001; // addi	$t0 $zero 65
		ram[66] = 32'B00011100000010000000000000000001; // sw	$t0 1($zero)
		ram[67] = 32'B00011000000101000000000000000000; // lw	$s0 0($zero)
		ram[68] = 32'B00011000000101010000000000000001; // lw	$s1 1($zero)
		ram[69] = 32'B00111110100101010100000000000000; // sbt	$t0 $s0 $s1
		ram[70] = 32'B00101001000000000000000000010000; // beq	$t0 0 L0
		ram[71] = 32'B00011000000101010000000000000000; // lw	$s1 0($zero)
		ram[72] = 32'B00011100000101010000000000000010; // sw	$s1 2($zero)
		ram[73] = 32'B00010100000000000000000000010011; // jump	L1
		ram[74] = 32'B00110000000000000000000000000000; // nop	L0
		ram[75] = 32'B00011000000101010000000000000001; // lw	$s1 1($zero)
		ram[76] = 32'B00011100000101010000000000000010; // sw	$s1 2($zero)
		ram[77] = 32'B00110000000000000000000000000000; // nop	L1
		ram[78] = 32'B00011000000101010000000000000010; // lw	$s1 2($zero)
		ram[79] = 32'B00001110101000100000000000000000; // move	$a0 $s1 
		ram[80] = 32'B00100100010000000000000000000000; // out	$a0  
		ram[81] = 32'B01110000000000000000000000000010; // Set PID 2	  
		ram[82] = 32'B01011000000000000000000000011000; // end file
		ram[83] = 32'B01010100000000000000000000000000; // begin file	  
		ram[84] = 32'B00001000000000010000000000000100; // addi	$ra $zero 4
		ram[85] = 32'B00001000000111110000000000011101; // addi	$sp $zero 29
		ram[86] = 32'B00010100000000000000000000000100; // jump	main
		ram[87] = 32'B00110000000000000000000000000000; // nop	main
		ram[88] = 32'B00001000000010000000000000000110; // addi	$t0 $zero 6
		ram[89] = 32'B00011100000010000000000000000001; // sw	$t0 1($zero)
		ram[90] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[91] = 32'B00011100000010000000000000000000; // sw	$t0 0($zero)
		ram[92] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[93] = 32'B00011100000010000000000000000010; // sw	$t0 2($zero)
		ram[94] = 32'B00110000000000000000000000000000; // nop	L0
		ram[95] = 32'B00011000000101000000000000000000; // lw	$s0 0($zero)
		ram[96] = 32'B00011000000101010000000000000001; // lw	$s1 1($zero)
		ram[97] = 32'B00010010100101010100000000000000; // slt	$t0 $s0 $s1
		ram[98] = 32'B00101001000000000000000000011110; // beq	$t0 0 L1
		ram[99] = 32'B00001000000010010000000000000010; // addi	$t1 $zero 2
		ram[100] = 32'B00011000000101010000000000000010; // lw	$s1 2($zero)
		ram[101] = 32'B00000001001101010101000000000010; // mult	$t2 $t1 $s1
		ram[102] = 32'B00011100000010100000000000000010; // sw	$t2 2($zero)
		ram[103] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[104] = 32'B00011000000101000000000000000000; // lw	$s0 0($zero)
		ram[105] = 32'B00000001000101000100100000000000; // add	$t1 $s0 $t0
		ram[106] = 32'B00011100000010010000000000000000; // sw	$t1 0($zero)
		ram[107] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[108] = 32'B00011000000101000000000000000010; // lw	$s0 2($zero)
		ram[109] = 32'B00000010100010000100100000000001; // sub	$t1 $s0 $t0
		ram[110] = 32'B00001101001000100000000000000000; // move	$a0 $t1 
		ram[111] = 32'B00100100010000000000000000000000; // out	$a0  
		ram[112] = 32'B00010100000000000000000000001011; // jump	L0
		ram[113] = 32'B00110000000000000000000000000000; // nop	L1
		ram[114] = 32'B00010100000000000000000000011111; // halt	  
		ram[115] = 32'B01011000000000000000000000110010; // end file	  		
		ram[116] = 32'B01100000000000000000000000000000; // HD_END
	end 

	always @ (posedge clk)
	begin
	
		// Write
		if (we)
			ram[addr] <= data;

		addr_reg <= addr;
	end
 
	assign q = ram[addr_reg];

endmodule
