module HDSimulado
#(parameter DATA_WIDTH=32, parameter ADDR_WIDTH=10)
(
	input [(DATA_WIDTH-1):0] data,
	input [(ADDR_WIDTH-1):0] addr,
	input we, clk,
	output [(DATA_WIDTH-1):0] q
);

	// Declare the RAM variable
	reg [DATA_WIDTH-1:0] ram[2**ADDR_WIDTH-1:0];

	// Variable to hold the registered read address
	reg [ADDR_WIDTH-1:0] addr_reg;

	initial 
	begin : INIT
		integer i;
		ram[ 0] = 32'B01010100000000000000000000000000; // begin file	  
		ram[ 1] = 32'B00001000000000010000000000011011; // addi	$ra $zero 27
		ram[ 2] = 32'B00001000000111110000000000110100; // addi	$sp $zero 52
		ram[ 3] = 32'B00010100000000000000000100010101; // jump	main
		ram[ 4] = 32'B00110000000000000000000000000000; // nop	Contexto
		ram[ 5] = 32'B00001000000111010000000111110100; // addi $z1, $zero, 500;
		ram[ 6] = 32'B00011111101000010000000000000000; // store $1,0($z1);
		ram[ 7] = 32'B00011111101000100000000000000001; // store $2,1($z1);
		ram[ 8] = 32'B00011111101000110000000000000010; // store $3,2($z1);
		ram[ 9] = 32'B00011111101001000000000000000011; // store $4,3($z1);
		ram[10] = 32'B00011111101001010000000000000100; // store $5,4($z1);
		ram[11] = 32'B00011111101001100000000000000101; // store $6,5($z1);
		ram[12] = 32'B00011111101001110000000000000110; // store $7,6($z1);
		ram[13] = 32'B00011111101010000000000000000111; // store $8,7($z1);
		ram[14] = 32'B00011111101010010000000000001000; // store $9,8($z1);
		ram[15] = 32'B00011111101010100000000000001001; // store $10,9($z1);
		ram[16] = 32'B00011111101010110000000000001010; // store $11,10($z1);
		ram[17] = 32'B00011111101011000000000000001011; // store $12,11($z1);
		ram[18] = 32'B00011111101011010000000000001100; // store $13,12($z1);
		ram[19] = 32'B00011111101011100000000000001101; // store $14,13($z1);
		ram[20] = 32'B00011111101011110000000000001110; // store $15,14($z1);
		ram[21] = 32'B00011111101100000000000000001111; // store $16,15($z1);
		ram[22] = 32'B00011111101100010000000000010000; // store $17,16($z1);
		ram[23] = 32'B00011111101100100000000000010001; // store $18,17($z1);
		ram[24] = 32'B00011111101100110000000000010010; // store $19,18($z1);
		ram[25] = 32'B00011111101101000000000000010011; // store $20,19($z1);
		ram[26] = 32'B00011111101101010000000000010100; // store $21,20($z1);
		ram[27] = 32'B00011111101101100000000000010101; // store $22,21($z1);
		ram[28] = 32'B00011111101101110000000000010110; // store $23,22($z1);
		ram[29] = 32'B00011111101110000000000000010111; // store $24,23($z1);
		ram[30] = 32'B00011111101110010000000000011000; // store $25,24($z1);
		ram[31] = 32'B00011111101110100000000000011001; // store $26,25($z1);
		ram[32] = 32'B00011111101110110000000000011010; // store $27,26($z1);
		ram[33] = 32'B00011111101111000000000000011011; // store $28,27($z1);
		ram[34] = 32'B00011111101111100000000000011100; // store $30,28($z1);
		ram[35] = 32'B00011111101111110000000000011110; // store $31,29($z1);
		ram[36] = 32'B00001000000111010000000000011111; // ADDI $z1,$zero,31
		ram[37] = 32'B00011000000111000000000000000010; // LOAD $z0,2($zero);
		ram[38] = 32'B00000011101111001110100000000010; // MULT $z1,$z1,$z0;
		ram[39] = 32'B00001011101111010000000111110100; // ADDI $z1,$z1,500
		ram[40] = 32'B00011011101000010000000000000000; // load $1,0($z1);
		ram[41] = 32'B00011011101000100000000000000001; // load $2,1($z1);
		ram[42] = 32'B00011011101000110000000000000010; // load $3,2($z1);
		ram[43] = 32'B00011011101001000000000000000011; // load $4,3($z1);
		ram[44] = 32'B00011011101001010000000000000100; // load $5,4($z1);
		ram[45] = 32'B00011011101001100000000000000101; // load $6,5($z1);
		ram[46] = 32'B00011011101001110000000000000110; // load $7,6($z1);
		ram[47] = 32'B00011011101010000000000000000111; // load $8,7($z1);
		ram[48] = 32'B00011011101010010000000000001000; // load $9,8($z1);
		ram[49] = 32'B00011011101010100000000000001001; // load $10,9($z1);
		ram[50] = 32'B00011011101010110000000000001010; // load $11,10($z1);
		ram[51] = 32'B00011011101011000000000000001011; // load $12,11($z1);
		ram[52] = 32'B00011011101011010000000000001100; // load $13,12($z1);
		ram[53] = 32'B00011011101011100000000000001101; // load $14,13($z1);
		ram[54] = 32'B00011011101011110000000000001110; // load $15,14($z1);
		ram[55] = 32'B00011011101100000000000000001111; // load $16,15($z1);
		ram[56] = 32'B00011011101100010000000000010000; // load $17,16($z1);
		ram[57] = 32'B00011011101100100000000000010001; // load $18,17($z1);
		ram[58] = 32'B00011011101100110000000000010010; // load $19,18($z1);
		ram[59] = 32'B00011011101101000000000000010011; // load $20,19($z1);
		ram[60] = 32'B00011011101101010000000000010100; // load $21,20($z1);
		ram[61] = 32'B00011011101101100000000000010101; // load $22,21($z1);
		ram[62] = 32'B00011011101101110000000000010110; // load $23,22($z1);
		ram[63] = 32'B00011011101110000000000000010111; // load $24,23($z1);
		ram[64] = 32'B00011011101110010000000000011000; // load $25,24($z1);
		ram[65] = 32'B00011011101110100000000000011001; // load $26,25($z1);
		ram[66] = 32'B00011011101110110000000000011010; // load $27,26($z1);
		ram[67] = 32'B00011011101111000000000000011011; // load $28,27($z1);
		ram[68] = 32'B00011011101111100000000000011100; // load $30,28($z1);
		ram[69] = 32'B00011011101111110000000000011101; // load $31,29($z1);
		ram[70] = 32'B00001000000111000000000000000001; // ADDI $z0,$zero,1;
		ram[71] = 32'B01110000000111000000000000000010; // SetPID $8 2($zero); -- Set_PID é um load na posicao alocada para ProcessoCorrente
		ram[72] = 32'B00011100000111000000000000000011;	// store $z0, $zero,3; 
		ram[73] = 32'B00001000000111010000000000011111; // ADDI $z1,$zero,31
		ram[74] = 32'B00011000000111000000000000000010; // LOAD $z0,2($zero);
		ram[75] = 32'B00000011101111001110100000000010; // MULT $z1,$z1,$z0;
		ram[76] = 32'B00001011101111010000000111110100; // ADDI $z1,$z1,500;
		ram[77] = 32'B00011111101000010000000000000000; // store $1,0($z1);
		ram[78] = 32'B00011111101000100000000000000001; // store $2,1($z1);
		ram[79] = 32'B00011111101000110000000000000010; // store $3,2($z1);
		ram[80] = 32'B00011111101001000000000000000011; // store $4,3($z1);
		ram[81] = 32'B00011111101001010000000000000100; // store $5,4($z1);
		ram[82] = 32'B00011111101001100000000000000101; // store $6,5($z1);
		ram[83] = 32'B00011111101001110000000000000110; // store $7,6($z1);
		ram[84] = 32'B00011111101010000000000000000111; // store $8,7($z1);
		ram[85] = 32'B00011111101010010000000000001000; // store $9,8($z1);
		ram[86] = 32'B00011111101010100000000000001001; // store $10,9($z1);
		ram[87] = 32'B00011111101010110000000000001010; // store $11,10($z1);
		ram[88] = 32'B00011111101011000000000000001011; // store $12,11($z1);
		ram[89] = 32'B00011111101011010000000000001100; // store $13,12($z1);
		ram[90] = 32'B00011111101011100000000000001101; // store $14,13($z1);
		ram[91] = 32'B00011111101011110000000000001110; // store $15,14($z1);
		ram[92] = 32'B00011111101100000000000000001111; // store $16,15($z1);
		ram[93] = 32'B00011111101100010000000000010000; // store $17,16($z1);
		ram[94] = 32'B00011111101100100000000000010001; // store $18,17($z1);
		ram[95] = 32'B00011111101100110000000000010010; // store $19,18($z1);
		ram[96] = 32'B00011111101101000000000000010011; // store $20,19($z1);
		ram[97] = 32'B00011111101101010000000000010100; // store $21,20($z1);
		ram[98] = 32'B00011111101101100000000000010101; // store $22,21($z1);
		ram[99] = 32'B00011111101101110000000000010110; // store $23,22($z1);
		ram[100] = 32'B00011111101110000000000000010111; // store $24,23($z1);
		ram[101] = 32'B00011111101110010000000000011000; // store $25,24($z1);
		ram[102] = 32'B00011111101110100000000000011001; // store $26,25($z1);
		ram[103] = 32'B00011111101110110000000000011010; // store $27,26($z1);
		ram[104] = 32'B00011111101111000000000000011011; // store $28,27($z1);
		ram[105] = 32'B00011111101111100000000000011100; // store $30,28($z1);
		ram[106] = 32'B00011111101111110000000000011101; // store $31,29($z1);
		ram[107] = 32'B00001000000111010000000111110100; // addi $z1, $zero, 500;
		ram[108] = 32'B00011011101000010000000000000000; // load $1,0($z1);
		ram[109] = 32'B00011011101000100000000000000001; // load $2,1($z1);
		ram[110] = 32'B00011011101000110000000000000010; // load $3,2($z1);
		ram[111] = 32'B00011011101001000000000000000011; // load $4,3($z1);
		ram[112] = 32'B00011011101001010000000000000100; // load $5,4($z1);
		ram[113] = 32'B00011011101001100000000000000101; // load $6,5($z1);
		ram[114] = 32'B00011011101001110000000000000110; // load $7,6($z1);
		ram[115] = 32'B00011011101010000000000000000111; // load $8,7($z1);
		ram[116] = 32'B00011011101010010000000000001000; // load $9,8($z1);
		ram[117] = 32'B00011011101010100000000000001001; // load $10,9($z1);
		ram[118] = 32'B00011011101010110000000000001010; // load $11,10($z1);
		ram[119] = 32'B00011011101011000000000000001011; // load $12,11($z1);
		ram[120] = 32'B00011011101011010000000000001100; // load $13,12($z1);
		ram[121] = 32'B00011011101011100000000000001101; // load $14,13($z1);
		ram[122] = 32'B00011011101011110000000000001110; // load $15,14($z1);
		ram[123] = 32'B00011011101100000000000000001111; // load $16,15($z1);
		ram[124] = 32'B00011011101100010000000000010000; // load $17,16($z1);
		ram[125] = 32'B00011011101100100000000000010001; // load $18,17($z1);
		ram[126] = 32'B00011011101100110000000000010010; // load $19,18($z1);
		ram[127] = 32'B00011011101101000000000000010011; // load $20,19($z1);
		ram[128] = 32'B00011011101101010000000000010100; // load $21,20($z1);
		ram[129] = 32'B00011011101101100000000000010101; // load $22,21($z1);
		ram[130] = 32'B00011011101101110000000000010110; // load $23,22($z1);
		ram[131] = 32'B00011011101110000000000000010111; // load $24,23($z1);
		ram[132] = 32'B00011011101110010000000000011000; // load $25,24($z1);
		ram[133] = 32'B00011011101110100000000000011001; // load $26,25($z1);
		ram[134] = 32'B00011011101110110000000000011010; // load $27,26($z1);
		ram[135] = 32'B00011011101111000000000000011011; // load $28,27($z1);
		ram[136] = 32'B00011011101111100000000000011100; // load $30,28($z1);
		ram[137] = 32'B00011011101111110000000000011110; // load $31,29($z1);  
		ram[138] = 32'B01010000001000010000000000000001; // subi	$ra $ra 1
		ram[139] = 32'B00011000001101000000000000000000; // lw	$s0 0($ra)
		ram[140] = 32'B01001110100000000000000000000000; // jr	$s0  
		ram[141] = 32'B00110000000000000000000000000000; // nop	InserirProcesso
		ram[142] = 32'B00011100000000100000000000001111; // sw	$a0 15($zero)
		ram[143] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[144] = 32'B00011000000101000000000000001111; // lw	$s0 15($zero)
		ram[145] = 32'B00000001000101000100100000000000; // add	$t1 $s0 $t0
		ram[146] = 32'B00011000000101010000000000000000; // lw	$s1 0($zero)
		ram[147] = 32'B00001010101010100000000000000100; // addi	$t2 $s1 4
		ram[148] = 32'B00011101010010010000000000000000; // sw	$t1 0($t2)
		ram[149] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[150] = 32'B00011000000101000000000000000000; // lw	$s0 0($zero)
		ram[151] = 32'B00000001000101000100100000000000; // add	$t1 $s0 $t0
		ram[152] = 32'B00011100000010010000000000000000; // sw	$t1 0($zero)
		ram[153] = 32'B01010000001000010000000000000001; // subi	$ra $ra 1
		ram[154] = 32'B00011000001101000000000000000000; // lw	$s0 0($ra)
		ram[155] = 32'B01001110100000000000000000000000; // jr	$s0  
		ram[156] = 32'B00110000000000000000000000000000; // nop	mod
		ram[157] = 32'B00011100000000100000000000010000; // sw	$a0 16($zero)
		ram[158] = 32'B00011100000000110000000000010001; // sw	$a1 17($zero)
		ram[159] = 32'B00011000000101000000000000010000; // lw	$s0 16($zero)
		ram[160] = 32'B00011000000101010000000000010001; // lw	$s1 17($zero)
		ram[161] = 32'B00000010100101010100000000000011; // div	$t0 $s0 $s1
		ram[162] = 32'B00011000000101010000000000010001; // lw	$s1 17($zero)
		ram[163] = 32'B00000001000101010100100000000010; // mult	$t1 $t0 $s1
		ram[164] = 32'B00011000000101000000000000010000; // lw	$s0 16($zero)
		ram[165] = 32'B00000010100010010101000000000001; // sub	$t2 $s0 $t1
		ram[166] = 32'B00001101010111100000000000000000; // move	$v0 $t2 
		ram[167] = 32'B01010000001000010000000000000001; // subi	$ra $ra 1
		ram[168] = 32'B00011000001101000000000000000000; // lw	$s0 0($ra)
		ram[169] = 32'B01001110100000000000000000000000; // jr	$s0  
		ram[170] = 32'B00110000000000000000000000000000; // nop	RoundRobinRun
		ram[171] = 32'B00001000000010110000000000000000; // addi	$t3 $zero 0
		ram[172] = 32'B00011100000010110000000000010010; // sw	$t3 18($zero)
		ram[173] = 32'B00110000000000000000000000000000; // nop	L0
		ram[174] = 32'B00001000000010000000000000000000; // addi	$t0 $zero 0
		ram[175] = 32'B00011000000101000000000000000000; // lw	$s0 0($zero)
		ram[176] = 32'B00111110100010000100100000000000; // sbt	$t1 $s0 $t0
		ram[177] = 32'B00101001001000000000000011100000; // beq	$t1 0 L1
		ram[178] = 32'B00011000000101010000000000010010; // lw	$s1 18($zero)
		ram[179] = 32'B00001110101000100000000000000000; // move	$a0 $s1 
		ram[180] = 32'B00011000000101010000000000000000; // lw	$s1 0($zero)
		ram[181] = 32'B00001110101000110000000000000000; // move	$a1 $s1 
		ram[182] = 32'B00001000000101000000000010111010; // addi	$s0 $zero 186
		ram[183] = 32'B00011100001101000000000000000000; // sw	$s0 0($ra)
		ram[184] = 32'B00001000001000010000000000000001; // addi	$ra $ra 1
		ram[185] = 32'B00010100000000000000000010011100; // jump	mod
		ram[186] = 32'B00011100000111100000000000010011; // sw	$v0 19($zero)
		ram[187] = 32'B00011000000101010000000000010011; // lw	$s1 19($zero)
		ram[188] = 32'B00011010101010000000000000000100; // lw	$t0 4($s1)
		ram[189] = 32'B00001000000010010000000000000000; // addi	$t1 $zero 0
		ram[190] = 32'B00111101000010010101000000000000; // sbt	$t2 $t0 $t1
		ram[191] = 32'B00101001010000000000000011011001; // beq	$t2 0 L2
		ram[192] = 32'B00011000000101010000000000010011; // lw	$s1 19($zero)
		ram[193] = 32'B00011010101010110000000000000100; // lw	$t3 4($s1)
		ram[194] = 32'B00011100000010110000000000000010; // sw	$t3 2($zero)
		ram[195] = 32'B00001000000101000000000011000111; // addi	$s0 $zero 199
		ram[196] = 32'B00011100001101000000000000000000; // sw	$s0 0($ra)
		ram[197] = 32'B00001000001000010000000000000001; // addi	$ra $ra 1
		ram[198] = 32'B00010100000000000000000000000100; // jump	Contexto
		ram[199] = 32'B00001000000010000000000000000000; // addi	$t0 $zero 0
		ram[200] = 32'B00011000000101000000000000000011; // lw	$s0 3($zero)
		ram[201] = 32'B01000010100010000100100000000000; // equal	$t1 $s0 $t0
		ram[202] = 32'B00101001001000000000000011010110; // beq	$t1 0 L4
		ram[203] = 32'B00001000000010100000000000000001; // addi	$t2 $zero 1
		ram[204] = 32'B00011100000010100000000000000011; // sw	$t2 3($zero)
		ram[205] = 32'B00011000000101010000000000010011; // lw	$s1 19($zero)
		ram[206] = 32'B00011010101010000000000000000100; // lw	$t0 4($s1)
		ram[207] = 32'B00001000000010010000000000000000; // addi	$t1 $zero 0
		ram[208] = 32'B01000001000010010101000000000000; // equal	$t2 $t0 $t1
		ram[209] = 32'B00001000000010110000000000000001; // addi	$t3 $zero 1
		ram[210] = 32'B00011000000101000000000000000000; // lw	$s0 0($zero)
		ram[211] = 32'B00000010100010110110000000000001; // sub	$t4 $s0 $t3
		ram[212] = 32'B00011100000011000000000000000000; // sw	$t4 0($zero)
		ram[213] = 32'B00010100000000000000000011010111; // jump	L5
		ram[214] = 32'B00110000000000000000000000000000; // nop	L4
		ram[215] = 32'B00110000000000000000000000000000; // nop	L5
		ram[216] = 32'B00010100000000000000000011011010; // jump	L3
		ram[217] = 32'B00110000000000000000000000000000; // nop	L2
		ram[218] = 32'B00110000000000000000000000000000; // nop	L3
		ram[219] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[220] = 32'B00011000000101000000000000010010; // lw	$s0 18($zero)
		ram[221] = 32'B00000001000101000100100000000000; // add	$t1 $s0 $t0
		ram[222] = 32'B00011100000010010000000000010010; // sw	$t1 18($zero)
		ram[223] = 32'B00010100000000000000000010101101; // jump	L0
		ram[224] = 32'B00110000000000000000000000000000; // nop	L1
		ram[225] = 32'B01010000001000010000000000000001; // subi	$ra $ra 1
		ram[226] = 32'B00011000001101000000000000000000; // lw	$s0 0($ra)
		ram[227] = 32'B01001110100000000000000000000000; // jr	$s0  
		ram[228] = 32'B00110000000000000000000000000000; // nop	SemPreempcao
		ram[229] = 32'B00001000000010000000000000000000; // addi	$t0 $zero 0
		ram[230] = 32'B00011100000010000000000000010110; // sw	$t0 22($zero)
		ram[231] = 32'B00110000000000000000000000000000; // nop	L6
		ram[232] = 32'B00001000000010000000000000000000; // addi	$t0 $zero 0
		ram[233] = 32'B00011000000101000000000000000000; // lw	$s0 0($zero)
		ram[234] = 32'B00111110100010000100100000000000; // sbt	$t1 $s0 $t0
		ram[235] = 32'B00101001001000000000000100010001; // beq	$t1 0 L7
		ram[236] = 32'B00110000000000000000000000000000; // nop	L8
		ram[237] = 32'B00011000000101010000000000010110; // lw	$s1 22($zero)
		ram[238] = 32'B00011010101010100000000000000100; // lw	$t2 4($s1)
		ram[239] = 32'B00001000000010110000000000000000; // addi	$t3 $zero 0
		ram[240] = 32'B00111101010010110110000000000000; // sbt	$t4 $t2 $t3
		ram[241] = 32'B00101001100000000000000100001011; // beq	$t4 0 L9
		ram[242] = 32'B00011000000101010000000000010110; // lw	$s1 22($zero)
		ram[243] = 32'B00011010101011010000000000000100; // lw	$t5 4($s1)
		ram[244] = 32'B00011100000011010000000000000010; // sw	$t5 2($zero)
		ram[245] = 32'B00001000000101000000000011111001; // addi	$s0 $zero 249
		ram[246] = 32'B00011100001101000000000000000000; // sw	$s0 0($ra)
		ram[247] = 32'B00001000001000010000000000000001; // addi	$ra $ra 1
		ram[248] = 32'B00010100000000000000000000000100; // jump	Contexto
		ram[249] = 32'B00001000000010000000000000000000; // addi	$t0 $zero 0
		ram[250] = 32'B00011000000101000000000000000011; // lw	$s0 3($zero)
		ram[251] = 32'B01000010100010000100100000000000; // equal	$t1 $s0 $t0
		ram[252] = 32'B00101001001000000000000100001000; // beq	$t1 0 L10
		ram[253] = 32'B00001000000010100000000000000001; // addi	$t2 $zero 1
		ram[254] = 32'B00011100000010100000000000000011; // sw	$t2 3($zero)
		ram[255] = 32'B00011000000101010000000000010110; // lw	$s1 22($zero)
		ram[256] = 32'B00011010101010000000000000000100; // lw	$t0 4($s1)
		ram[257] = 32'B00001000000010010000000000000000; // addi	$t1 $zero 0
		ram[258] = 32'B01000001000010010101000000000000; // equal	$t2 $t0 $t1
		ram[259] = 32'B00001000000010110000000000000001; // addi	$t3 $zero 1
		ram[260] = 32'B00011000000101000000000000000000; // lw	$s0 0($zero)
		ram[261] = 32'B00000010100010110110000000000001; // sub	$t4 $s0 $t3
		ram[262] = 32'B00011100000011000000000000000000; // sw	$t4 0($zero)
		ram[263] = 32'B00010100000000000000000100001001; // jump	L11
		ram[264] = 32'B00110000000000000000000000000000; // nop	L10
		ram[265] = 32'B00110000000000000000000000000000; // nop	L11
		ram[266] = 32'B00010100000000000000000011101100; // jump	L8
		ram[267] = 32'B00110000000000000000000000000000; // nop	L9
		ram[268] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[269] = 32'B00011000000101000000000000010110; // lw	$s0 22($zero)
		ram[270] = 32'B00000001000101000100100000000000; // add	$t1 $s0 $t0
		ram[271] = 32'B00011100000010010000000000010110; // sw	$t1 22($zero)
		ram[272] = 32'B00010100000000000000000011100111; // jump	L6
		ram[273] = 32'B00110000000000000000000000000000; // nop	L7
		ram[274] = 32'B01010000001000010000000000000001; // subi	$ra $ra 1
		ram[275] = 32'B00011000001101000000000000000000; // lw	$s0 0($ra)
		ram[276] = 32'B01001110100000000000000000000000; // jr	$s0  
		ram[277] = 32'B00110000000000000000000000000000; // nop	main
		ram[278] = 32'B00001000000010000000000000000000; // addi	$t0 $zero 0
		ram[279] = 32'B00011100000010000000000000000000; // sw	$t0 0($zero)
		ram[280] = 32'B00001000000010000000000000000000; // addi	$t0 $zero 0
		ram[281] = 32'B00011100000010000000000000011000; // sw	$t0 24($zero)
		ram[282] = 32'B00011000000101010000000000011000; // lw	$s1 24($zero)
		ram[283] = 32'B00001110101000100000000000000000; // move	$a0 $s1 
		ram[284] = 32'B00001000000101000000000100100000; // addi	$s0 $zero 288
		ram[285] = 32'B00011100001101000000000000000000; // sw	$s0 0($ra)
		ram[286] = 32'B00001000001000010000000000000001; // addi	$ra $ra 1
		ram[287] = 32'B00010100000000000000000010001101; // jump	InserirProcesso
		ram[288] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[289] = 32'B00011100000010000000000000011000; // sw	$t0 24($zero)
		ram[290] = 32'B00011000000101010000000000011000; // lw	$s1 24($zero)
		ram[291] = 32'B00001110101000100000000000000000; // move	$a0 $s1 
		ram[292] = 32'B00001000000101000000000100101000; // addi	$s0 $zero 296
		ram[293] = 32'B00011100001101000000000000000000; // sw	$s0 0($ra)
		ram[294] = 32'B00001000001000010000000000000001; // addi	$ra $ra 1
		ram[295] = 32'B00010100000000000000000010001101; // jump	InserirProcesso
		ram[296] = 32'B00001000000010000000000000000010; // addi	$t0 $zero 2
		ram[297] = 32'B00011100000010000000000000011000; // sw	$t0 24($zero)
		ram[298] = 32'B00011000000101010000000000011000; // lw	$s1 24($zero)
		ram[299] = 32'B00001110101000100000000000000000; // move	$a0 $s1 
		ram[300] = 32'B00001000000101000000000100110000; // addi	$s0 $zero 304
		ram[301] = 32'B00011100001101000000000000000000; // sw	$s0 0($ra)
		ram[302] = 32'B00001000001000010000000000000001; // addi	$ra $ra 1
		ram[303] = 32'B00010100000000000000000010001101; // jump	InserirProcesso
		ram[304] = 32'B00001000000101000000000100110100; // addi	$s0 $zero 308
		ram[305] = 32'B00011100001101000000000000000000; // sw	$s0 0($ra)
		ram[306] = 32'B00001000001000010000000000000001; // addi	$ra $ra 1
		ram[307] = 32'B00010100000000000000000010101010; // jump	RoundRobinRun
		ram[308] = 32'B00110000000000000000000000000000; // nop	L12
		ram[309] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[310] = 32'B00001000000010010000000000000001; // addi	$t1 $zero 1
		ram[311] = 32'B01000001000010010101000000000000; // equal	$t2 $t0 $t1
		ram[312] = 32'B00101001010000000000000100111010; // beq	$t2 0 L13
		ram[313] = 32'B00010100000000000000000100110100; // jump	L12
		ram[314] = 32'B00110000000000000000000000000000; // nop	L13
		ram[315] = 32'B00001000000111010000000000000001; // addi	$s9 $zero 1
		ram[316] = 32'B10000100000111000000000000000000; // move	$s8 $zero 
		ram[317] = 32'B01011000000000000000000000110010; // end file	  
		ram[318] = 32'B00110000000000000000000000000000;
		ram[319] = 32'B00110000000000000000000000000000;
		ram[320] = 32'B00110000000000000000000000000000;
		ram[321] = 32'B01010100000000000000000000000000; // begin file	  
		ram[322] = 32'B00001000000000010000000000001000; // addi	$ra $zero 8
		ram[323] = 32'B00001000000111110000000000100001; // addi	$sp $zero 33
		ram[324] = 32'B00010100000000000000000000101001; // jump	main
		ram[325] = 32'B00110000000000000000000000000000; // nop	Combinatoria
		ram[326] = 32'B00011100000000100000000000000000; // sw	$a0 0($zero)
		ram[327] = 32'B00011100000000110000000000000001; // sw	$a1 1($zero)
		ram[328] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[329] = 32'B00011100000010000000000000000010; // sw	$t0 2($zero)
		ram[330] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[331] = 32'B00011100000010000000000000000011; // sw	$t0 3($zero)
		ram[332] = 32'B00110000000000000000000000000000; // nop	L0
		ram[333] = 32'B00001000000010000000000000000000; // addi	$t0 $zero 0
		ram[334] = 32'B00011000000101000000000000000001; // lw	$s0 1($zero)
		ram[335] = 32'B00111110100010000100100000000000; // sbt	$t1 $s0 $t0
		ram[336] = 32'B00101001001000000000000000100001; // beq	$t1 0 L1
		ram[337] = 32'B00011000000101000000000000000010; // lw	$s0 2($zero)
		ram[338] = 32'B00011000000101010000000000000000; // lw	$s1 0($zero)
		ram[339] = 32'B00000010100101010101000000000010; // mult	$t2 $s0 $s1
		ram[340] = 32'B00011100000010100000000000000010; // sw	$t2 2($zero)
		ram[341] = 32'B00011000000101000000000000000011; // lw	$s0 3($zero)
		ram[342] = 32'B00011000000101010000000000000001; // lw	$s1 1($zero)
		ram[343] = 32'B00000010100101010100000000000010; // mult	$t0 $s0 $s1
		ram[344] = 32'B00011100000010000000000000000011; // sw	$t0 3($zero)
		ram[345] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[346] = 32'B00011000000101000000000000000000; // lw	$s0 0($zero)
		ram[347] = 32'B00000010100010000100100000000001; // sub	$t1 $s0 $t0
		ram[348] = 32'B00011100000010010000000000000000; // sw	$t1 0($zero)
		ram[349] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[350] = 32'B00011000000101000000000000000001; // lw	$s0 1($zero)
		ram[351] = 32'B00000010100010000100100000000001; // sub	$t1 $s0 $t0
		ram[352] = 32'B00011100000010010000000000000001; // sw	$t1 1($zero)
		ram[353] = 32'B00010100000000000000000000001011; // jump	L0
		ram[354] = 32'B00110000000000000000000000000000; // nop	L1
		ram[355] = 32'B00011000000101000000000000000010; // lw	$s0 2($zero)
		ram[356] = 32'B00011000000101010000000000000011; // lw	$s1 3($zero)
		ram[357] = 32'B00000010100101010100000000000011; // div	$t0 $s0 $s1
		ram[358] = 32'B00001101000111100000000000000000; // move	$v0 $t0 
		ram[359] = 32'B01010000001000010000000000000001; // subi	$ra $ra 1
		ram[360] = 32'B00011000001101000000000000000000; // lw	$s0 0($ra)
		ram[361] = 32'B01001110100000000000000000000000; // jr	$s0  
		ram[362] = 32'B00110000000000000000000000000000; // nop	main
		ram[363] = 32'B00001000000010010000000000001111; // addi	$t1 $zero 15
		ram[364] = 32'B00011100000010010000000000000100; // sw	$t1 4($zero)
		ram[365] = 32'B00001000000010000000000000000110; // addi	$t0 $zero 6
		ram[366] = 32'B00011100000010000000000000000101; // sw	$t0 5($zero)
		ram[367] = 32'B00011000000101010000000000000100; // lw	$s1 4($zero)
		ram[368] = 32'B00001110101000100000000000000000; // move	$a0 $s1 
		ram[369] = 32'B00011000000101010000000000000101; // lw	$s1 5($zero)
		ram[370] = 32'B00001110101000110000000000000000; // move	$a1 $s1 
		ram[371] = 32'B00001000000101000000000000110110; // addi	$s0 $zero 54
		ram[372] = 32'B00011100001101000000000000000000; // sw	$s0 0($ra)
		ram[373] = 32'B00001000001000010000000000000001; // addi	$ra $ra 1
		ram[374] = 32'B00010100000000000000000000000100; // jump	Combinatoria
		ram[375] = 32'B00001111110001000000000000000000; // move	$a2 $v0 
		ram[376] = 32'B00100100100000000000000000000000; // out	$a2  
		ram[377] = 32'B00001000000111010000000000000001; // addi	$s9 $zero 1
		ram[378] = 32'B10000100000111000000000000000000; // kernel_swap	  
		ram[379] = 32'B01011000000000000000000000110010; // end file	 
		ram[380] = 32'B01010100000000000000000000000000; // begin file	  
		ram[381] = 32'B00001000000000010000000000000101; // addi	$ra $zero 5
		ram[382] = 32'B00001000000111110000000000011110; // addi	$sp $zero 30
		ram[383] = 32'B00010100000000000000000000000100; // jump	main
		ram[384] = 32'B00110000000000000000000000000000; // nop	main
		ram[385] = 32'B00001000000010000000000000000010; // addi	$t0 $zero 2
		ram[386] = 32'B00011100000010000000000000000000; // sw	$t0 0($zero)
		ram[387] = 32'B00001000000010000000000000000111; // addi	$t0 $zero 7
		ram[388] = 32'B00011100000010000000000000000001; // sw	$t0 1($zero)
		ram[389] = 32'B00011000000101010000000000000001; // lw	$s1 1($zero)
		ram[390] = 32'B00011100000101010000000000000010; // sw	$s1 2($zero)
		ram[391] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[392] = 32'B00011100000010000000000000000011; // sw	$t0 3($zero)
		ram[393] = 32'B00110000000000000000000000000000; // nop	L0
		ram[394] = 32'B00001000000010000000000000000000; // addi	$t0 $zero 0
		ram[395] = 32'B00011000000101000000000000000010; // lw	$s0 2($zero)
		ram[396] = 32'B00111110100010000100100000000000; // sbt	$t1 $s0 $t0
		ram[397] = 32'B00101001001000000000000000011011; // beq	$t1 0 L1
		ram[398] = 32'B00011000000101000000000000000011; // lw	$s0 3($zero)
		ram[399] = 32'B00011000000101010000000000000000; // lw	$s1 0($zero)
		ram[400] = 32'B00000010100101010101000000000010; // mult	$t2 $s0 $s1
		ram[401] = 32'B00011100000010100000000000000011; // sw	$t2 3($zero)
		ram[402] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[403] = 32'B00011000000101000000000000000010; // lw	$s0 2($zero)
		ram[404] = 32'B00000010100010000100100000000001; // sub	$t1 $s0 $t0
		ram[405] = 32'B00011100000010010000000000000010; // sw	$t1 2($zero)
		ram[406] = 32'B00010100000000000000000000001101; // jump	L0
		ram[407] = 32'B00110000000000000000000000000000; // nop	L1
		ram[408] = 32'B00011000000101010000000000000011; // lw	$s1 3($zero)
		ram[409] = 32'B00001110101000100000000000000000; // move	$a0 $s1 
		ram[410] = 32'B00100100010000000000000000000000; // out	$a0  
		ram[411] = 32'B00001000000111010000000000000001; // addi	$s9 $zero 1
		ram[412] = 32'B10000100000111000000000000000000; // kernel_swap	  
		ram[413] = 32'B01011000000000000000000000110010; // end file	 
		ram[414] = 32'B01010100000000000000000000000000; // begin file	  
		ram[415] = 32'B00001000000000010000000000000100; // addi	$ra $zero 4
		ram[416] = 32'B00001000000111110000000000011101; // addi	$sp $zero 29
		ram[417] = 32'B00010100000000000000000000000100; // jump	main
		ram[418] = 32'B00110000000000000000000000000000; // nop	main
		ram[419] = 32'B00001000000010000000000000000110; // addi	$t0 $zero 6
		ram[420] = 32'B00011100000010000000000000000001; // sw	$t0 1($zero)
		ram[421] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[422] = 32'B00011100000010000000000000000000; // sw	$t0 0($zero)
		ram[423] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[424] = 32'B00011100000010000000000000000010; // sw	$t0 2($zero)
		ram[425] = 32'B00110000000000000000000000000000; // nop	L0
		ram[426] = 32'B00011000000101000000000000000000; // lw	$s0 0($zero)
		ram[427] = 32'B00011000000101010000000000000001; // lw	$s1 1($zero)
		ram[428] = 32'B00010010100101010100000000000000; // slt	$t0 $s0 $s1
		ram[429] = 32'B00101001000000000000000000011110; // beq	$t0 0 L1
		ram[430] = 32'B00001000000010010000000000000010; // addi	$t1 $zero 2
		ram[431] = 32'B00011000000101010000000000000010; // lw	$s1 2($zero)
		ram[432] = 32'B00000001001101010101000000000010; // mult	$t2 $t1 $s1
		ram[433] = 32'B00011100000010100000000000000010; // sw	$t2 2($zero)
		ram[434] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[435] = 32'B00011000000101000000000000000000; // lw	$s0 0($zero)
		ram[436] = 32'B00000001000101000100100000000000; // add	$t1 $s0 $t0
		ram[437] = 32'B00011100000010010000000000000000; // sw	$t1 0($zero)
		ram[438] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		ram[439] = 32'B00011000000101000000000000000010; // lw	$s0 2($zero)
		ram[440] = 32'B00000010100010000100100000000001; // sub	$t1 $s0 $t0
		ram[441] = 32'B00001101001000100000000000000000; // move	$a0 $t1 
		ram[442] = 32'B00100100010000000000000000000000; // out	$a0  
		ram[443] = 32'B00010100000000000000000000001011; // jump	L0
		ram[444] = 32'B00110000000000000000000000000000; // nop	L1
		ram[445] = 32'B00001000000111010000000000000001; // addi	$s9 $zero 1
		ram[446] = 32'B10000100000111000000000000000000; // kernel_swap	  
		ram[447] = 32'B01011000000000000000000000110010; // end file	  
		ram[448] = 32'B01100000000000000000000000000000; // HD_END
	end 

	always @ (posedge clk)
	begin
	
		// Write
		if (we)
			ram[addr] <= data;

		addr_reg <= addr;
	end
 
	assign q = ram[addr_reg];

endmodule
